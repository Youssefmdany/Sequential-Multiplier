module adder(input[15:0] dataa,datab,output[15:0] sum);



assign sum = dataa + datab;

endmodule 